class packet;

    randc bit [3:0]a;
	randc bit [3:0]b;
	
	bit y1,y2,y3;
	
	/* bit [3:0]prev_a,prev_b;
	
	constraint c1{a!=prev_a;b!=prev_b;}
	
	
	function void post_randomize();
	a=prev_a;
	b=prev_b;
	endfunction */
	
	
	
	
	endclass
